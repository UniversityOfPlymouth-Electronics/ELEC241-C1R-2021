library ieee;
use ieee.std_logic_1164.all;

entity mux21 is


	port 
	(
		SEL   : in std_logic;
		A0		: in std_logic;
		A1    : in std_logic;

		Q   	: out std_logic
	);

end entity;

architecture rtl of mux21 is

begin

	-- write code here
	
end rtl;
